magic
tech scmos
timestamp 1770733275
<< nwell >>
rect -14 -17 16 9
<< polysilicon >>
rect -3 -4 -1 -2
rect 1 -4 3 -2
rect -3 -34 -1 -12
rect 1 -19 3 -12
rect 1 -23 2 -19
rect 6 -23 7 -19
rect 5 -34 7 -23
rect -3 -40 -1 -38
rect 5 -40 7 -38
<< ndiffusion >>
rect -4 -38 -3 -34
rect -1 -38 0 -34
rect 4 -38 5 -34
rect 7 -38 8 -34
<< pdiffusion >>
rect -5 -12 -3 -4
rect -1 -12 1 -4
rect 3 -12 5 -4
rect 9 -12 13 -4
<< metal1 >>
rect -14 6 16 9
rect -14 2 -9 6
rect -5 2 0 6
rect 4 2 8 6
rect 12 2 16 6
rect -14 -1 16 2
rect -9 -4 -5 -1
rect 4 -12 5 -4
rect -14 -23 2 -19
rect 9 -26 13 -4
rect -14 -30 -7 -26
rect 0 -31 13 -26
rect 0 -34 4 -31
rect -8 -41 -4 -38
rect 8 -41 12 -38
rect -12 -43 16 -41
rect -12 -47 -8 -43
rect -4 -47 0 -43
rect 4 -47 8 -43
rect 12 -47 16 -43
rect -12 -56 16 -47
<< ntransistor >>
rect -3 -38 -1 -34
rect 5 -38 7 -34
<< ptransistor >>
rect -3 -12 -1 -4
rect 1 -12 3 -4
<< polycontact >>
rect -7 -30 -3 -26
rect 2 -23 6 -19
<< ndcontact >>
rect -8 -38 -4 -34
rect 0 -38 4 -34
rect 8 -38 12 -34
<< pdcontact >>
rect -9 -12 -5 -4
rect 5 -12 9 -4
<< psubstratepcontact >>
rect -8 -47 -4 -43
rect 0 -47 4 -43
rect 8 -47 12 -43
<< nsubstratencontact >>
rect -9 2 -5 6
rect 0 2 4 6
rect 8 2 12 6
<< labels >>
rlabel metal1 13 3 13 3 7 VDD
rlabel metal1 11 -24 11 -24 7 out
rlabel metal1 -13 -21 -13 -21 3 A
rlabel metal1 -12 -28 -12 -28 3 B
rlabel metal1 14 -46 14 -46 7 GND
<< end >>
