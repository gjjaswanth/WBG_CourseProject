magic
tech scmos
timestamp 1770742332
<< nwell >>
rect -3 -4 36 9
<< polysilicon >>
rect 9 7 12 11
rect 21 7 24 11
rect 9 -20 12 -1
rect 21 -20 24 -1
rect 9 -32 12 -28
rect 21 -32 24 -28
<< ndiffusion >>
rect 1 -22 9 -20
rect 1 -26 3 -22
rect 7 -26 9 -22
rect 1 -28 9 -26
rect 12 -28 21 -20
rect 24 -23 34 -20
rect 24 -28 27 -23
rect 32 -28 34 -23
<< pdiffusion >>
rect 0 5 9 7
rect 0 1 3 5
rect 7 1 9 5
rect 0 -1 9 1
rect 12 5 21 7
rect 12 0 14 5
rect 19 0 21 5
rect 12 -1 21 0
rect 24 5 32 7
rect 24 1 27 5
rect 31 1 32 5
rect 24 -1 32 1
<< metal1 >>
rect 3 17 31 18
rect 7 13 14 17
rect 18 13 25 17
rect 29 13 31 17
rect 3 12 31 13
rect 3 5 7 12
rect 27 5 31 12
rect 14 -10 19 0
rect 14 -15 32 -10
rect 3 -35 7 -26
rect 27 -23 32 -15
rect 3 -36 36 -35
rect 3 -40 4 -36
rect 8 -40 13 -36
rect 17 -40 21 -36
rect 25 -40 29 -36
rect 33 -40 36 -36
rect 3 -41 36 -40
<< ntransistor >>
rect 9 -28 12 -20
rect 21 -28 24 -20
<< ptransistor >>
rect 9 -1 12 7
rect 21 -1 24 7
<< ndcontact >>
rect 3 -26 7 -22
rect 27 -28 32 -23
<< pdcontact >>
rect 3 1 7 5
rect 14 0 19 5
rect 27 1 31 5
<< psubstratepcontact >>
rect 4 -40 8 -36
rect 13 -40 17 -36
rect 21 -40 25 -36
rect 29 -40 33 -36
<< nsubstratencontact >>
rect 3 13 7 17
rect 14 13 18 17
rect 25 13 29 17
<< end >>
