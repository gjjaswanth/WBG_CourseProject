* SPICE3 file created from nand3.ext - technology: scmos

.model pfet pmos level=1 VTO=-0.7 KP=40u LAMBDA=0.02
.model nfet nmos level=1 VTO=0.7 KP=80u LAMBDA=0.02
.option scale=1u

*======================
* Transistors (corrected nodes and bulks)

M1000 out A vdd vdd pfet w=8 l=3
+  ad=36p pd=17u as=72p ps=34u

M1003 out B vdd vdd pfet w=8 l=3
+  ad=64p pd=32u as=36p ps=17u

M1001 out B a_12_n28# 0 nfet w=8 l=3
+  ad=80p pd=36u as=36p ps=17u

M1002 a_12_n28# A 0 0 nfet w=8 l=3
+  ad=36p pd=17u as=64p ps=32u


*======================
* Power Supply
VDD_SRC vdd 0 5

* Input A
VA A 0 PULSE(0 5 0n 1n 1n 20n 40n)

* Input B
VB B 0 PULSE(0 5 0n 1n 1n 40n 80n)

* Output load
CL out 0 10f

*======================
* Analysis
.tran 1n 200n

.control
run
plot V(A)
plot V(B)
plot V(out)
.endc

.end

