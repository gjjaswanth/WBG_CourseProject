magic
tech scmos
timestamp 1770524022
<< nwell >>
rect -10 4 11 27
<< polysilicon >>
rect -2 14 0 16
rect -2 1 0 6
rect -1 -3 0 1
rect -2 -9 0 -3
rect -2 -16 0 -13
<< ndiffusion >>
rect -3 -13 -2 -9
rect 0 -13 3 -9
rect 7 -13 8 -9
<< pdiffusion >>
rect -7 13 -2 14
rect -3 9 -2 13
rect -7 6 -2 9
rect 0 12 8 14
rect 0 8 3 12
rect 7 8 8 12
rect 0 6 8 8
<< metal1 >>
rect -10 21 -7 25
rect -3 21 1 25
rect 5 21 7 25
rect -10 20 7 21
rect -7 13 -3 20
rect 3 1 7 8
rect -10 -3 -5 1
rect 3 -3 12 1
rect 3 -9 7 -3
rect -7 -18 -3 -13
rect -3 -22 2 -18
rect 6 -22 7 -18
<< ntransistor >>
rect -2 -13 0 -9
<< ptransistor >>
rect -2 6 0 14
<< polycontact >>
rect -5 -3 -1 1
<< ndcontact >>
rect -7 -13 -3 -9
rect 3 -13 7 -9
<< pdcontact >>
rect -7 9 -3 13
rect 3 8 7 12
<< psubstratepcontact >>
rect -7 -22 -3 -18
rect 2 -22 6 -18
<< nsubstratencontact >>
rect -7 21 -3 25
rect 1 21 5 25
<< labels >>
rlabel metal1 -1 -20 -1 -20 1 gnd!
rlabel metal1 -1 22 -1 22 5 vdd!
rlabel metal1 -10 -3 -10 1 3 in
rlabel metal1 12 -3 12 1 7 out
<< end >>
